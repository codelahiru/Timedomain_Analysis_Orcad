** Profile: "SCHEMATIC1-biaspoint_sim2"  [ F:\Projects\Orcad Capture CIS\Project_0005\Timedomain_Analysis_Orcad\Time_Domain_Analysis-PSpiceFiles\SCHEMATIC1\biaspoint_sim2.sim ] 

** Creating circuit file "biaspoint_sim2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Gayan Lahiru\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
